module nor_gate(O,A,B);
  input A,B;
  output O;
  nor(O,A,B);
endmodule