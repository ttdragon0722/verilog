module nand_gate(O,A,B);
  input A,B;
  output O;
  nand(O,A,B);
endmodule